module test_mod01_bonus;

tester tester();

endmodule

