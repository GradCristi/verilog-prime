module test_add_10;

tester tester();

endmodule

