module test_call_bonus;

tester tester();

endmodule

