module test_add_immediate;

tester tester();

endmodule

