module test_jcond;

tester tester();

endmodule

