module test_jmp_10;

tester tester();

endmodule

