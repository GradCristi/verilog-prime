module test_jmp_simple_00;

tester tester();

endmodule

