module test_jmp_simple_11;

tester tester();

endmodule

