module test_jcond_simple;

tester tester();

endmodule

