module test_inc_10;

tester tester();

endmodule

