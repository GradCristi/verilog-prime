module test_push_10;

tester tester();

endmodule

