module test_mov_immediate;

tester tester();

endmodule

