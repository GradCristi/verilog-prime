module test_mov_10;

tester tester();

endmodule

