module test_pf_bonus;

tester tester();

endmodule

