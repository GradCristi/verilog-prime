module test_push_simple;

tester tester();

endmodule

