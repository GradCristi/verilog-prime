module test_mov_simple;

tester tester();

endmodule

